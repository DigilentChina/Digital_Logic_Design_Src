module gates4a_tb;
  reg [3:0] a;
  wire [5:0] y;
  gates4a uut(a,y);
  initial
    begin
      a = 4'b0000; #100;
      a = 4'b0001; #100;
      a = 4'b0010; #100;
      a = 4'b0011; #100;
      a = 4'b0100; #100;
      a = 4'b0101; #100;
      a = 4'b0110; #100;
      a = 4'b0111; #100;
      a = 4'b1000; #100;
      a = 4'b1001; #100;
      a = 4'b1010; #100;
      a = 4'b1011; #100;
      a = 4'b1100; #100;
      a = 4'b1101; #100;
      a = 4'b1110; #100;
      a = 4'b1111;
    end
endmodule